netcdf parameters { // parameters file in CDL

dimensions:

variables:
  int scenario_id;
  int NX, NY, NZ;
  double hX, hY, hZ, V, ir_const;
  double vw, vo, swc, sor;
  int St, Pt, ND;
  int solver_inner, solver_outer;

data:
  scenario_id = 1;

  NX = 10;

  NY = 10;

  NZ = 2;

  hX = 6.096000000;

  hY = 3.048000000;

  hZ = 0.609600000;

  V = 0.1132673863680000e2;

  ir_const = 0.7085561497326203e-3;

  vw = 3e-4;

  vo = 3e-3;

  swc = 0.2000;

  sor = 0.2000;

  St = 5;

  Pt = 100;

  ND = 2000;

  solver_inner = 64;

  solver_outer = 100000;

}